package parameters is

  constant dmem_size : integer := 1024;

  constant code_bin_path : string := "code.bin";

end package parameters;
